module test_aryan;
    reg [1:0] in1, in2, in3;
    wire [1:0] out;
    wire error;

    voter voter_instance (in1, in2, in3, out, error);

    initial begin
        in1 = 2'd0;    in2 = 2'd0;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd0;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd0;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd0;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd1;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd1;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd1;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd1;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd2;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd2;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd2;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd2;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd3;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd3;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd3;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd0;    in2 = 2'd3;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd0;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd0;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd0;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd0;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd1;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd1;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd1;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd1;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd2;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd2;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd2;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd2;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd3;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd3;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd3;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd1;    in2 = 2'd3;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd0;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd0;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd0;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd0;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd1;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd1;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd1;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd1;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd2;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd2;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd2;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd2;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd3;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd3;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd3;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd2;    in2 = 2'd3;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd0;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd0;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd0;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd0;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd1;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd1;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd1;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd1;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd2;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd2;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd2;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd2;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd3;    in3 = 2'd0;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd3;    in3 = 2'd1;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd3;    in3 = 2'd2;
        #1 $display("%b %b", out, error);
        in1 = 2'd3;    in2 = 2'd3;    in3 = 2'd3;
        #1 $display("%b %b", out, error);
    end
endmodule
