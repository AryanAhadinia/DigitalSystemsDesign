module test;
    reg     [31:0]  data;
    reg             data_ready;
    reg             clk;
    reg             reset;
    reg     [31:0]  constant;
    reg     [3:0]   opcode;

    wire    [31:0]  out;
    wire    out_valid;

    procesor    pcs (data, data_ready, clk, reset, constant, opcode, out, out_valid);

    initial begin
        clk = 1'b0;
    end
    always begin
        #5 clk = !clk;
    end

    initial begin
        // ADD
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b0010;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;

        #10	data = 32'b01101111110001000000001111000011;
        #10	data = 32'b10010011110010111001111010001111;
        #10	data = 32'b11010100001110110100101001100011;
        #10	data = 32'b11101010001010011111101011101001;
        #10	data = 32'b10101000110000000111100111100001;
        #10	data = 32'b10011000111010000110001111000010;
        #10	data = 32'b00100101110010110011001011111001;
        #10	data = 32'b00101001000101010000100001001011;
        #100

        // SUB
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b0011;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;

        #10	data = 32'b01101111110001000000001111000011;
        #10	data = 32'b10010011110010111001111010001111;
        #10	data = 32'b11010100001110110100101001100011;
        #10	data = 32'b11101010001010011111101011101001;
        #10	data = 32'b10101000110000000111100111100001;
        #10	data = 32'b10011000111010000110001111000010;
        #10	data = 32'b00100101110010110011001011111001;
        #10	data = 32'b00101001000101010000100001001011;
        #100

        // MUL
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b0001;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;

        #10	data = 32'b01101111110001000000001111000011;
        #10	data = 32'b10010011110010111001111010001111;
        #10	data = 32'b11010100001110110100101001100011;
        #10	data = 32'b11101010001010011111101011101001;
        #10	data = 32'b10101000110000000111100111100001;
        #10	data = 32'b10011000111010000110001111000010;
        #10	data = 32'b00100101110010110011001011111001;
        #10	data = 32'b00101001000101010000100001001011;
        #100

        // AND
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b1101;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;

        #10	data = 32'b01101111110001000000001111000011;
        #10	data = 32'b10010011110010111001111010001111;
        #10	data = 32'b11010100001110110100101001100011;
        #10	data = 32'b11101010001010011111101011101001;
        #10	data = 32'b10101000110000000111100111100001;
        #10	data = 32'b10011000111010000110001111000010;
        #10	data = 32'b00100101110010110011001011111001;
        #10	data = 32'b00101001000101010000100001001011;
        #100

        // XOR
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b1111;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;

        #10	data = 32'b01101111110001000000001111000011;
        #10	data = 32'b10010011110010111001111010001111;
        #10	data = 32'b11010100001110110100101001100011;
        #10	data = 32'b11101010001010011111101011101001;
        #10	data = 32'b10101000110000000111100111100001;
        #10	data = 32'b10011000111010000110001111000010;
        #10	data = 32'b00100101110010110011001011111001;
        #10	data = 32'b00101001000101010000100001001011;
        #100

        // SDC
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b1000;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;
        #100

        // SRR
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b1001;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;
        #100

        // SUC
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b1010;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;
        #100

        // SLR
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b1011;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;
        #100

        // NOP
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        data_ready = 1'b1;
        opcode = 4'b0000;
        #100

        // AWC
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        constant = 32'b11010101101011100100000101111011;
        data_ready = 1'b1;
        opcode = 4'b1100;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;
        #100

        // XWC
        #1  reset = 1'b1;
        #1  reset = 1'b0;
        constant = 32'b11010101101011100100000101111011;
        data_ready = 1'b1;
        opcode = 4'b1110;
        #3	data = 32'b11010101101011100100000101111011;
        #10	data = 32'b10111001010011110011110001100011;
        #10	data = 32'b11110001001111100100011001110001;
        #10	data = 32'b11000000111100110100000111101101;
        #10	data = 32'b01000110110100010000001000000000;
        #10	data = 32'b11001010011100001001101010101000;
        #10	data = 32'b10110010011010111001011101111110;
        #10	data = 32'b11001010111111011110010100000001;
        #100

        $stop;

    end

    always @(posedge out_valid) begin
        $display("Begin");
        #10 $display("%b", out);
        #10 $display("%b", out);
        #10 $display("%b", out);
        #10 $display("%b", out);
        #10 $display("%b", out);
        #10 $display("%b", out);
        #10 $display("%b", out);
        #10 $display("%b", out);
        $display("End");
    end
endmodule
