module test_aryan;
    wire [7:0] m;
    reg [3:0] a;
    reg [3:0] b;

    unsigned_multiplier ump (m, a, b);

    initial begin
        $monitor($time, "\t%d = %d * %d", m, a, b);
        #1  a = 4'd0;   b = 4'd0;
        #1  a = 4'd0;   b = 4'd1;
        #1  a = 4'd0;   b = 4'd2;
        #1  a = 4'd0;   b = 4'd3;
        #1  a = 4'd0;   b = 4'd4;
        #1  a = 4'd0;   b = 4'd5;
        #1  a = 4'd0;   b = 4'd6;
        #1  a = 4'd0;   b = 4'd7;
        #1  a = 4'd0;   b = 4'd8;
        #1  a = 4'd0;   b = 4'd9;
        #1  a = 4'd0;   b = 4'd10;
        #1  a = 4'd0;   b = 4'd11;
        #1  a = 4'd0;   b = 4'd12;
        #1  a = 4'd0;   b = 4'd13;
        #1  a = 4'd0;   b = 4'd14;
        #1  a = 4'd0;   b = 4'd15;
        #1  a = 4'd1;   b = 4'd0;
        #1  a = 4'd1;   b = 4'd1;
        #1  a = 4'd1;   b = 4'd2;
        #1  a = 4'd1;   b = 4'd3;
        #1  a = 4'd1;   b = 4'd4;
        #1  a = 4'd1;   b = 4'd5;
        #1  a = 4'd1;   b = 4'd6;
        #1  a = 4'd1;   b = 4'd7;
        #1  a = 4'd1;   b = 4'd8;
        #1  a = 4'd1;   b = 4'd9;
        #1  a = 4'd1;   b = 4'd10;
        #1  a = 4'd1;   b = 4'd11;
        #1  a = 4'd1;   b = 4'd12;
        #1  a = 4'd1;   b = 4'd13;
        #1  a = 4'd1;   b = 4'd14;
        #1  a = 4'd1;   b = 4'd15;
        #1  a = 4'd2;   b = 4'd0;
        #1  a = 4'd2;   b = 4'd1;
        #1  a = 4'd2;   b = 4'd2;
        #1  a = 4'd2;   b = 4'd3;
        #1  a = 4'd2;   b = 4'd4;
        #1  a = 4'd2;   b = 4'd5;
        #1  a = 4'd2;   b = 4'd6;
        #1  a = 4'd2;   b = 4'd7;
        #1  a = 4'd2;   b = 4'd8;
        #1  a = 4'd2;   b = 4'd9;
        #1  a = 4'd2;   b = 4'd10;
        #1  a = 4'd2;   b = 4'd11;
        #1  a = 4'd2;   b = 4'd12;
        #1  a = 4'd2;   b = 4'd13;
        #1  a = 4'd2;   b = 4'd14;
        #1  a = 4'd2;   b = 4'd15;
        #1  a = 4'd3;   b = 4'd0;
        #1  a = 4'd3;   b = 4'd1;
        #1  a = 4'd3;   b = 4'd2;
        #1  a = 4'd3;   b = 4'd3;
        #1  a = 4'd3;   b = 4'd4;
        #1  a = 4'd3;   b = 4'd5;
        #1  a = 4'd3;   b = 4'd6;
        #1  a = 4'd3;   b = 4'd7;
        #1  a = 4'd3;   b = 4'd8;
        #1  a = 4'd3;   b = 4'd9;
        #1  a = 4'd3;   b = 4'd10;
        #1  a = 4'd3;   b = 4'd11;
        #1  a = 4'd3;   b = 4'd12;
        #1  a = 4'd3;   b = 4'd13;
        #1  a = 4'd3;   b = 4'd14;
        #1  a = 4'd3;   b = 4'd15;
        #1  a = 4'd4;   b = 4'd0;
        #1  a = 4'd4;   b = 4'd1;
        #1  a = 4'd4;   b = 4'd2;
        #1  a = 4'd4;   b = 4'd3;
        #1  a = 4'd4;   b = 4'd4;
        #1  a = 4'd4;   b = 4'd5;
        #1  a = 4'd4;   b = 4'd6;
        #1  a = 4'd4;   b = 4'd7;
        #1  a = 4'd4;   b = 4'd8;
        #1  a = 4'd4;   b = 4'd9;
        #1  a = 4'd4;   b = 4'd10;
        #1  a = 4'd4;   b = 4'd11;
        #1  a = 4'd4;   b = 4'd12;
        #1  a = 4'd4;   b = 4'd13;
        #1  a = 4'd4;   b = 4'd14;
        #1  a = 4'd4;   b = 4'd15;
        #1  a = 4'd5;   b = 4'd0;
        #1  a = 4'd5;   b = 4'd1;
        #1  a = 4'd5;   b = 4'd2;
        #1  a = 4'd5;   b = 4'd3;
        #1  a = 4'd5;   b = 4'd4;
        #1  a = 4'd5;   b = 4'd5;
        #1  a = 4'd5;   b = 4'd6;
        #1  a = 4'd5;   b = 4'd7;
        #1  a = 4'd5;   b = 4'd8;
        #1  a = 4'd5;   b = 4'd9;
        #1  a = 4'd5;   b = 4'd10;
        #1  a = 4'd5;   b = 4'd11;
        #1  a = 4'd5;   b = 4'd12;
        #1  a = 4'd5;   b = 4'd13;
        #1  a = 4'd5;   b = 4'd14;
        #1  a = 4'd5;   b = 4'd15;
        #1  a = 4'd6;   b = 4'd0;
        #1  a = 4'd6;   b = 4'd1;
        #1  a = 4'd6;   b = 4'd2;
        #1  a = 4'd6;   b = 4'd3;
        #1  a = 4'd6;   b = 4'd4;
        #1  a = 4'd6;   b = 4'd5;
        #1  a = 4'd6;   b = 4'd6;
        #1  a = 4'd6;   b = 4'd7;
        #1  a = 4'd6;   b = 4'd8;
        #1  a = 4'd6;   b = 4'd9;
        #1  a = 4'd6;   b = 4'd10;
        #1  a = 4'd6;   b = 4'd11;
        #1  a = 4'd6;   b = 4'd12;
        #1  a = 4'd6;   b = 4'd13;
        #1  a = 4'd6;   b = 4'd14;
        #1  a = 4'd6;   b = 4'd15;
        #1  a = 4'd7;   b = 4'd0;
        #1  a = 4'd7;   b = 4'd1;
        #1  a = 4'd7;   b = 4'd2;
        #1  a = 4'd7;   b = 4'd3;
        #1  a = 4'd7;   b = 4'd4;
        #1  a = 4'd7;   b = 4'd5;
        #1  a = 4'd7;   b = 4'd6;
        #1  a = 4'd7;   b = 4'd7;
        #1  a = 4'd7;   b = 4'd8;
        #1  a = 4'd7;   b = 4'd9;
        #1  a = 4'd7;   b = 4'd10;
        #1  a = 4'd7;   b = 4'd11;
        #1  a = 4'd7;   b = 4'd12;
        #1  a = 4'd7;   b = 4'd13;
        #1  a = 4'd7;   b = 4'd14;
        #1  a = 4'd7;   b = 4'd15;
        #1  a = 4'd8;   b = 4'd0;
        #1  a = 4'd8;   b = 4'd1;
        #1  a = 4'd8;   b = 4'd2;
        #1  a = 4'd8;   b = 4'd3;
        #1  a = 4'd8;   b = 4'd4;
        #1  a = 4'd8;   b = 4'd5;
        #1  a = 4'd8;   b = 4'd6;
        #1  a = 4'd8;   b = 4'd7;
        #1  a = 4'd8;   b = 4'd8;
        #1  a = 4'd8;   b = 4'd9;
        #1  a = 4'd8;   b = 4'd10;
        #1  a = 4'd8;   b = 4'd11;
        #1  a = 4'd8;   b = 4'd12;
        #1  a = 4'd8;   b = 4'd13;
        #1  a = 4'd8;   b = 4'd14;
        #1  a = 4'd8;   b = 4'd15;
        #1  a = 4'd9;   b = 4'd0;
        #1  a = 4'd9;   b = 4'd1;
        #1  a = 4'd9;   b = 4'd2;
        #1  a = 4'd9;   b = 4'd3;
        #1  a = 4'd9;   b = 4'd4;
        #1  a = 4'd9;   b = 4'd5;
        #1  a = 4'd9;   b = 4'd6;
        #1  a = 4'd9;   b = 4'd7;
        #1  a = 4'd9;   b = 4'd8;
        #1  a = 4'd9;   b = 4'd9;
        #1  a = 4'd9;   b = 4'd10;
        #1  a = 4'd9;   b = 4'd11;
        #1  a = 4'd9;   b = 4'd12;
        #1  a = 4'd9;   b = 4'd13;
        #1  a = 4'd9;   b = 4'd14;
        #1  a = 4'd9;   b = 4'd15;
        #1  a = 4'd10;   b = 4'd0;
        #1  a = 4'd10;   b = 4'd1;
        #1  a = 4'd10;   b = 4'd2;
        #1  a = 4'd10;   b = 4'd3;
        #1  a = 4'd10;   b = 4'd4;
        #1  a = 4'd10;   b = 4'd5;
        #1  a = 4'd10;   b = 4'd6;
        #1  a = 4'd10;   b = 4'd7;
        #1  a = 4'd10;   b = 4'd8;
        #1  a = 4'd10;   b = 4'd9;
        #1  a = 4'd10;   b = 4'd10;
        #1  a = 4'd10;   b = 4'd11;
        #1  a = 4'd10;   b = 4'd12;
        #1  a = 4'd10;   b = 4'd13;
        #1  a = 4'd10;   b = 4'd14;
        #1  a = 4'd10;   b = 4'd15;
        #1  a = 4'd11;   b = 4'd0;
        #1  a = 4'd11;   b = 4'd1;
        #1  a = 4'd11;   b = 4'd2;
        #1  a = 4'd11;   b = 4'd3;
        #1  a = 4'd11;   b = 4'd4;
        #1  a = 4'd11;   b = 4'd5;
        #1  a = 4'd11;   b = 4'd6;
        #1  a = 4'd11;   b = 4'd7;
        #1  a = 4'd11;   b = 4'd8;
        #1  a = 4'd11;   b = 4'd9;
        #1  a = 4'd11;   b = 4'd10;
        #1  a = 4'd11;   b = 4'd11;
        #1  a = 4'd11;   b = 4'd12;
        #1  a = 4'd11;   b = 4'd13;
        #1  a = 4'd11;   b = 4'd14;
        #1  a = 4'd11;   b = 4'd15;
        #1  a = 4'd12;   b = 4'd0;
        #1  a = 4'd12;   b = 4'd1;
        #1  a = 4'd12;   b = 4'd2;
        #1  a = 4'd12;   b = 4'd3;
        #1  a = 4'd12;   b = 4'd4;
        #1  a = 4'd12;   b = 4'd5;
        #1  a = 4'd12;   b = 4'd6;
        #1  a = 4'd12;   b = 4'd7;
        #1  a = 4'd12;   b = 4'd8;
        #1  a = 4'd12;   b = 4'd9;
        #1  a = 4'd12;   b = 4'd10;
        #1  a = 4'd12;   b = 4'd11;
        #1  a = 4'd12;   b = 4'd12;
        #1  a = 4'd12;   b = 4'd13;
        #1  a = 4'd12;   b = 4'd14;
        #1  a = 4'd12;   b = 4'd15;
        #1  a = 4'd13;   b = 4'd0;
        #1  a = 4'd13;   b = 4'd1;
        #1  a = 4'd13;   b = 4'd2;
        #1  a = 4'd13;   b = 4'd3;
        #1  a = 4'd13;   b = 4'd4;
        #1  a = 4'd13;   b = 4'd5;
        #1  a = 4'd13;   b = 4'd6;
        #1  a = 4'd13;   b = 4'd7;
        #1  a = 4'd13;   b = 4'd8;
        #1  a = 4'd13;   b = 4'd9;
        #1  a = 4'd13;   b = 4'd10;
        #1  a = 4'd13;   b = 4'd11;
        #1  a = 4'd13;   b = 4'd12;
        #1  a = 4'd13;   b = 4'd13;
        #1  a = 4'd13;   b = 4'd14;
        #1  a = 4'd13;   b = 4'd15;
        #1  a = 4'd14;   b = 4'd0;
        #1  a = 4'd14;   b = 4'd1;
        #1  a = 4'd14;   b = 4'd2;
        #1  a = 4'd14;   b = 4'd3;
        #1  a = 4'd14;   b = 4'd4;
        #1  a = 4'd14;   b = 4'd5;
        #1  a = 4'd14;   b = 4'd6;
        #1  a = 4'd14;   b = 4'd7;
        #1  a = 4'd14;   b = 4'd8;
        #1  a = 4'd14;   b = 4'd9;
        #1  a = 4'd14;   b = 4'd10;
        #1  a = 4'd14;   b = 4'd11;
        #1  a = 4'd14;   b = 4'd12;
        #1  a = 4'd14;   b = 4'd13;
        #1  a = 4'd14;   b = 4'd14;
        #1  a = 4'd14;   b = 4'd15;
        #1  a = 4'd15;   b = 4'd0;
        #1  a = 4'd15;   b = 4'd1;
        #1  a = 4'd15;   b = 4'd2;
        #1  a = 4'd15;   b = 4'd3;
        #1  a = 4'd15;   b = 4'd4;
        #1  a = 4'd15;   b = 4'd5;
        #1  a = 4'd15;   b = 4'd6;
        #1  a = 4'd15;   b = 4'd7;
        #1  a = 4'd15;   b = 4'd8;
        #1  a = 4'd15;   b = 4'd9;
        #1  a = 4'd15;   b = 4'd10;
        #1  a = 4'd15;   b = 4'd11;
        #1  a = 4'd15;   b = 4'd12;
        #1  a = 4'd15;   b = 4'd13;
        #1  a = 4'd15;   b = 4'd14;
        #1  a = 4'd15;   b = 4'd15;
    end  
endmodule
